module day_05

pub fn solve_first(input string) string {
	return input
}

pub fn solve_second(input string) string {
	return input
}
